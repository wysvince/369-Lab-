`timescale 1ns / 1ps

module HDU();

endmodule;